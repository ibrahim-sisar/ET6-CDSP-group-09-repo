measure,Country,cause,metric,year,Deaths Val,upper,lower
Deaths,China,COVID-19,Percent,2021,9.170442215509476e-05,0.0003320497854356,7.303893605064585e-06
Deaths,China,COVID-19,Rate,2021,0.0747041830796572,0.2828000127164385,0.0060046003698948
Deaths,Italy,COVID-19,Percent,2021,0.0908639792683596,0.0956988571689352,0.0865860908207042
Deaths,Italy,COVID-19,Rate,2021,106.19180038529572,111.9663099106196,100.9876724355437
Deaths,Chile,COVID-19,Percent,2021,0.2091465729864521,0.2177875615323765,0.1997087082862726
Deaths,Chile,COVID-19,Rate,2021,149.0404092460287,154.8478180973691,143.25717266713886
Deaths,Japan,COVID-19,Percent,2021,0.0103558601051742,0.0123227147925933,0.0087398157575816
Deaths,Japan,COVID-19,Rate,2021,11.657724081474315,13.872192365649909,9.849034458573955
Deaths,United States of America,COVID-19,Percent,2021,0.1392929867018255,0.1424576424126143,0.1365513067551055
Deaths,United States of America,COVID-19,Rate,2021,145.35398147932767,148.75147847625857,142.6152141492136
Deaths,Nigeria,COVID-19,Percent,2021,0.0718631535545515,0.0833613832137604,0.0612248779422539
Deaths,Nigeria,COVID-19,Rate,2021,56.44638552029111,63.663965276931336,50.52948134269381
Deaths,India,COVID-19,Percent,2021,0.1420160570163332,0.1530028210195809,0.1311158724472252
Deaths,India,COVID-19,Rate,2021,117.80370068827496,122.76382986126136,111.8438189725278
Deaths,Egypt,COVID-19,Percent,2021,0.1551880366822783,0.2049674857334592,0.1015254759787769
Deaths,Egypt,COVID-19,Rate,2021,103.96988609236828,134.62148530750758,68.96838754624139
Deaths,Italy,COVID-19,Percent,2020,0.1130485348610423,0.1170980158214756,0.1089868815583398
Deaths,Italy,COVID-19,Rate,2020,139.2720837898269,144.3082847151729,134.12932973358335
Deaths,Japan,COVID-19,Percent,2020,0.0025412593754785,0.0028706142677613,0.0022726000789291
Deaths,Japan,COVID-19,Rate,2020,2.71456126331636,3.0703090618549123,2.423480203519094
Deaths,China,COVID-19,Percent,2020,0.0023674046023309,0.0117635580402405,0.0005064345390425
Deaths,China,COVID-19,Rate,2020,1.8988807796412688,9.668453975892492,0.4137580881263417
Deaths,Nigeria,COVID-19,Percent,2020,0.0493641058280502,0.0559062024319146,0.0421641479808037
Deaths,Nigeria,COVID-19,Rate,2020,38.63730895990837,42.25435843765667,35.625862475744206
Deaths,Chile,COVID-19,Percent,2020,0.1694455223097943,0.1770027522243449,0.1619435510756737
Deaths,Chile,COVID-19,Rate,2020,112.95868489361132,118.06204026503823,108.00838610174942
Deaths,United States of America,COVID-19,Percent,2020,0.1270171103227867,0.1315621711807492,0.1225722281896749
Deaths,United States of America,COVID-19,Rate,2020,128.64146045427427,133.47057198116588,124.07161118760182
Deaths,India,COVID-19,Percent,2020,0.0903649591715642,0.0977827916046732,0.0821034459208865
Deaths,India,COVID-19,Rate,2020,68.6771185506763,72.66079819100513,64.50467827413775
Deaths,Egypt,COVID-19,Percent,2020,0.1100951012091408,0.1448001749234581,0.0741228321084871
Deaths,Egypt,COVID-19,Rate,2020,68.19287875990663,90.14021015607231,47.07465288102832
